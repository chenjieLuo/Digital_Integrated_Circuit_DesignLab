
module chenjie_module_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n4;
  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  ENI U2 ( .A(carry[7]), .B(n4), .Z(SUM[7]) );
  IVI U1 ( .A(A[7]), .Z(n4) );
  IVI U3 ( .A(A[0]), .Z(SUM[0]) );
endmodule


module chenjie_module_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  IVI U2 ( .A(n12), .Z(n1) );
  IVI U3 ( .A(n1), .Z(n2) );
  IVDA U4 ( .A(A[6]), .Z(n3) );
  IVI U5 ( .A(A[0]), .Z(n5) );
  IVI U6 ( .A(n5), .Z(n6) );
  IVI U7 ( .A(A[0]), .Z(n7) );
  IVI U8 ( .A(n6), .Z(SUM[0]) );
  ENI U9 ( .A(n8), .B(A[7]), .Z(SUM[7]) );
  ND2I U10 ( .A(n9), .B(n10), .Z(n8) );
  NR2I U11 ( .A(n25), .B(n11), .Z(n10) );
  ND2I U12 ( .A(A[3]), .B(A[2]), .Z(n11) );
  NR2I U13 ( .A(n12), .B(n13), .Z(n9) );
  ND2I U14 ( .A(A[5]), .B(A[6]), .Z(n13) );
  ENI U15 ( .A(n14), .B(n3), .Z(SUM[6]) );
  ND2I U16 ( .A(n15), .B(n16), .Z(n14) );
  NR2I U17 ( .A(n7), .B(n17), .Z(n16) );
  ND2I U18 ( .A(A[1]), .B(A[2]), .Z(n17) );
  NR2I U19 ( .A(n18), .B(n19), .Z(n15) );
  ND2I U20 ( .A(A[4]), .B(A[5]), .Z(n19) );
  ENI U21 ( .A(A[5]), .B(n20), .Z(SUM[5]) );
  ND2I U22 ( .A(n21), .B(n22), .Z(n20) );
  NR2I U23 ( .A(n5), .B(n23), .Z(n22) );
  ND2I U24 ( .A(A[4]), .B(A[3]), .Z(n23) );
  AN2I U25 ( .A(A[1]), .B(A[2]), .Z(n21) );
  ENI U26 ( .A(n24), .B(n2), .Z(SUM[4]) );
  IVI U27 ( .A(A[4]), .Z(n12) );
  NR2I U28 ( .A(n28), .B(n11), .Z(n24) );
  ND2I U29 ( .A(A[1]), .B(A[0]), .Z(n25) );
  ENI U30 ( .A(n26), .B(n18), .Z(SUM[3]) );
  IVI U31 ( .A(A[3]), .Z(n18) );
  NR2I U32 ( .A(n7), .B(n27), .Z(n26) );
  ND2I U33 ( .A(A[1]), .B(A[2]), .Z(n27) );
  ENI U34 ( .A(A[2]), .B(n28), .Z(SUM[2]) );
  ND2I U35 ( .A(A[1]), .B(A[0]), .Z(n28) );
  ENI U36 ( .A(n6), .B(n29), .Z(SUM[1]) );
  IVI U37 ( .A(A[1]), .Z(n29) );
endmodule


module chenjie_module ( clk, reset, throttle, set, accel, coast, cancel, 
        resume, brake, speed, cruise_speed, cruise_on );
  output [7:0] speed;
  output [7:0] cruise_speed;
  input clk, reset, throttle, set, accel, coast, cancel, resume, brake;
  output cruise_on;
  wire   n838, n2669, n839, n840, n841, n842, n843, n844, n845, N36, N37, N38,
         N39, N40, N41, N42, N43, N46, N47, N48, N49, N50, N51, N52, N53, N197,
         N198, N200, N201, N202, N255, N257, N259, N261, N263, N267, n159,
         n166, n168, n169, n170, n174, n176, n178, n179, n180, n1231, n1307,
         n1311, n1474, n1738, n1852, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2068, n2069, n2070, n2072, n2073, n2075, n2076, n2077, n2078, n2079,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668;
  assign speed[4] = n838;
  assign cruise_speed[5] = n840;
  assign cruise_speed[4] = n841;
  assign cruise_speed[2] = n843;
  assign cruise_speed[1] = n844;
  assign cruise_speed[0] = n845;

  FD1 \cached_speed_reg[0]  ( .D(n2661), .CP(set), .Q(n2027) );
  FD1 cruise_on_reg ( .D(n2228), .CP(clk), .Q(cruise_on) );
  FD1 \speed_reg[7]  ( .D(n180), .CP(clk), .Q(speed[7]), .QN(n2240) );
  FD1 \speed_reg[6]  ( .D(n179), .CP(clk), .Q(speed[6]), .QN(n2268) );
  FD1 \cruise_speed_reg[0]  ( .D(n2111), .CP(clk), .Q(n845), .QN(n2262) );
  FD1 \cruise_speed_reg[7]  ( .D(n2662), .CP(clk), .Q(cruise_speed[7]), .QN(
        n159) );
  FD1 \speed_reg[5]  ( .D(n178), .CP(clk), .Q(speed[5]) );
  FD1 \speed_reg[4]  ( .D(n1738), .CP(clk), .Q(n838), .QN(n2028) );
  FD1 \speed_reg[3]  ( .D(n176), .CP(clk), .Q(speed[3]) );
  FD1 \speed_reg[0]  ( .D(n2663), .CP(clk), .Q(speed[0]) );
  FD1 \speed_reg[1]  ( .D(n174), .CP(clk), .Q(speed[1]), .QN(n2072) );
  FD1 \speed_reg[2]  ( .D(n1311), .CP(clk), .Q(n2669), .QN(n2073) );
  FD1 \cached_speed_reg[1]  ( .D(n2664), .CP(set), .Q(n2023), .QN(n2089) );
  FD1 \cached_speed_reg[2]  ( .D(n2665), .CP(set), .Q(n2022) );
  FD1 \cached_speed_reg[3]  ( .D(n170), .CP(set), .Q(n2021) );
  FD1 \cached_speed_reg[4]  ( .D(n169), .CP(set), .Q(n2020), .QN(n2090) );
  FD1 \cached_speed_reg[5]  ( .D(n168), .CP(set), .Q(n2024) );
  FD1 \cached_speed_reg[6]  ( .D(n2666), .CP(set), .Q(n2025) );
  FD1 \cruise_speed_reg[6]  ( .D(n2098), .CP(clk), .Q(n839), .QN(n2140) );
  FD1 \cruise_speed_reg[5]  ( .D(n2099), .CP(clk), .Q(n840), .QN(n2137) );
  FD1 \cruise_speed_reg[1]  ( .D(n2041), .CP(clk), .Q(n844), .QN(n2265) );
  FD1 \cruise_speed_reg[2]  ( .D(n2039), .CP(clk), .Q(n843), .QN(n2266) );
  FD1 \cruise_speed_reg[3]  ( .D(n2040), .CP(clk), .Q(n842), .QN(n2086) );
  FD1 \cruise_speed_reg[4]  ( .D(n2038), .CP(clk), .Q(n841), .QN(n2019) );
  FD1 \cached_speed_reg[7]  ( .D(n166), .CP(set), .Q(n2026), .QN(n2091) );
  chenjie_module_DW01_inc_0 r97 ( .A({n2029, n1474, n2030, n2031, n2250, n2668, 
        n2168, n2032}), .SUM({N43, N42, N41, N40, N39, N38, N37, N36}) );
  chenjie_module_DW01_inc_1 add_43 ( .A({N255, N257, N259, N261, N263, n2260, 
        N267, n2263}), .SUM({N53, N52, N51, N50, N49, N48, N47, N46}) );
  INVX4 U815 ( .A(n2060), .Y(n2055) );
  NAND2X1 U816 ( .A(n2247), .B(n2397), .Y(n2033) );
  ND2I U817 ( .A(n2605), .B(n2037), .Z(n2034) );
  ND2I U818 ( .A(n2034), .B(n2035), .Z(n2171) );
  OR2P U819 ( .A(n2036), .B(n2634), .Z(n2035) );
  IVI U820 ( .A(n2094), .Z(n2036) );
  AN2I U821 ( .A(n2606), .B(n2094), .Z(n2037) );
  MUX21LP U822 ( .A(n2609), .B(n2608), .S(brake), .Z(n2611) );
  ND2I U823 ( .A(n2526), .B(n2525), .Z(n2038) );
  OR2X2 U824 ( .A(n2399), .B(n2400), .Y(n2185) );
  ND2I U825 ( .A(n2542), .B(n2541), .Z(n2039) );
  ND2I U826 ( .A(n2534), .B(n2533), .Z(n2040) );
  ND2I U827 ( .A(n2548), .B(n2547), .Z(n2041) );
  IVDA U828 ( .A(n2361), .Y(n2042), .Z(n2043) );
  IVDA U829 ( .A(n2354), .Y(n2044), .Z(n2045) );
  IVDA U830 ( .A(N47), .Y(n2046), .Z(n2047) );
  OR2I U831 ( .A(n2109), .B(n2046), .Z(n2048) );
  B2IP U832 ( .A(n2365), .Z2(n2049) );
  B4IP U833 ( .A(n2368), .Z(n2051) );
  B2I U834 ( .A(n2144), .Z1(n2052), .Z2(n2053) );
  AN2I U835 ( .A(n2446), .B(n2495), .Z(n2054) );
  BUFX2 U836 ( .A(n2403), .Y(n2056) );
  NAND3X1 U837 ( .A(n2208), .B(n2209), .C(n2055), .Y(n2057) );
  MUX21L U838 ( .A(speed[5]), .B(N41), .S(n2121), .Z(n2413) );
  AN2I U839 ( .A(resume), .B(n2188), .Z(n2058) );
  NAND2X1 U840 ( .A(n2244), .B(n2212), .Y(n2059) );
  AND2X2 U841 ( .A(n2113), .B(n2404), .Y(n2060) );
  NAND2X1 U842 ( .A(n2033), .B(n2063), .Y(n2061) );
  AND2X1 U843 ( .A(n2185), .B(n2401), .Y(n2062) );
  AND2X1 U844 ( .A(n2185), .B(n2402), .Y(n2063) );
  B4I U845 ( .A(n2142), .Z(n2144) );
  AND2X1 U846 ( .A(n2110), .B(n2056), .Y(n2114) );
  B5IP U847 ( .A(n2232), .Z(n2395) );
  B5IP U848 ( .A(n2229), .Z(n2402) );
  ND2I U849 ( .A(n2065), .B(n2079), .Z(n2229) );
  B5IP U850 ( .A(n2222), .Z(n2404) );
  ND2I U851 ( .A(n2078), .B(n2223), .Z(n2222) );
  IVI U852 ( .A(n2369), .Z(n2370) );
  IVI U853 ( .A(n2644), .Z(n2093) );
  AO7 U854 ( .A(n1852), .B(n2597), .C(speed[5]), .Z(n2269) );
  AN2I U855 ( .A(n2451), .B(n2450), .Z(n2064) );
  OR2I U856 ( .A(n2515), .B(n2109), .Z(n2065) );
  B2I U857 ( .A(n842), .Z2(cruise_speed[3]) );
  B2I U858 ( .A(n2614), .Z1(n2068), .Z2(n2069) );
  B2IP U859 ( .A(n2367), .Z2(n2070) );
  B2IP U860 ( .A(n2406), .Z2(n2220) );
  AN2I U861 ( .A(n2456), .B(n2156), .Z(n2075) );
  AN2I U862 ( .A(n2470), .B(n2469), .Z(n2076) );
  IVDA U863 ( .A(n2390), .Y(n2077) );
  OR2I U864 ( .A(n2129), .B(n2140), .Z(n2078) );
  AN2I U865 ( .A(n2380), .B(n2379), .Z(n2079) );
  B2I U866 ( .A(n839), .Z2(cruise_speed[6]) );
  IVDA U867 ( .A(N53), .Y(n2082), .Z(n2083) );
  IVDA U868 ( .A(N52), .Y(n2084), .Z(n2085) );
  AN2I U869 ( .A(n2500), .B(n2499), .Z(n2087) );
  AN2I U870 ( .A(n2466), .B(n2465), .Z(n2088) );
  IVI U871 ( .A(accel), .Z(n2145) );
  ND2I U872 ( .A(n2106), .B(n2092), .Z(n2126) );
  NR2I U873 ( .A(n2097), .B(n2646), .Z(n2092) );
  ENI U874 ( .A(n2647), .B(n2093), .Z(n2639) );
  AN2I U875 ( .A(n2635), .B(n2196), .Z(n2094) );
  MUX21LP U876 ( .A(n2064), .B(n2097), .S(brake), .Z(n2237) );
  ND2I U877 ( .A(n2514), .B(n2117), .Z(n2095) );
  OR2I U878 ( .A(n2096), .B(n2582), .Z(n2489) );
  ND2I U879 ( .A(n2479), .B(n2483), .Z(n2096) );
  ND2I U880 ( .A(n2105), .B(n2602), .Z(n2097) );
  IVI U881 ( .A(n2132), .Z(n2103) );
  ND2I U882 ( .A(n2565), .B(n2564), .Z(n2098) );
  ND2I U883 ( .A(n2557), .B(n2556), .Z(n2099) );
  ND2I U884 ( .A(n2511), .B(n2656), .Z(n2100) );
  OR2I U885 ( .A(n2138), .B(n2172), .Z(n2101) );
  OR2I U886 ( .A(n2138), .B(n2578), .Z(n2102) );
  AN2I U887 ( .A(n2103), .B(n2104), .Z(n2105) );
  NR2I U888 ( .A(n2138), .B(n2578), .Z(n2104) );
  ND2I U889 ( .A(n2106), .B(n2605), .Z(n2647) );
  NR2I U890 ( .A(n2604), .B(n2637), .Z(n2106) );
  AND2X1 U891 ( .A(n2360), .B(n2030), .Y(n2217) );
  ND2I U892 ( .A(n2381), .B(n2344), .Z(n2107) );
  IVI U893 ( .A(n2107), .Z(n2267) );
  BUFX2 U894 ( .A(n2369), .Y(n2108) );
  IVI U895 ( .A(n2177), .Z(n2273) );
  MUX21LP U896 ( .A(N47), .B(n844), .S(n2145), .Z(n2278) );
  IVI U897 ( .A(n2133), .Z(n2109) );
  MUX21LP U898 ( .A(n2277), .B(n2276), .S(accel), .Z(n2279) );
  IVAP U899 ( .A(n2377), .Z(n2110) );
  ND2I U900 ( .A(n2359), .B(n2358), .Z(n2377) );
  MUX21LP U901 ( .A(N51), .B(n840), .S(n2145), .Z(n2297) );
  ND2I U902 ( .A(n2632), .B(n2631), .Z(n2111) );
  ND2I U903 ( .A(coast), .B(n2284), .Z(n2112) );
  NAND2X1 U904 ( .A(n2243), .B(n2059), .Y(n2113) );
  IVI U905 ( .A(n2130), .Z(n2115) );
  ND2I U906 ( .A(coast), .B(n2127), .Z(n2116) );
  ND2I U907 ( .A(set), .B(n2510), .Z(n2117) );
  IVAP U908 ( .A(n2195), .Z(n2410) );
  AN2I U909 ( .A(n842), .B(n2518), .Z(N263) );
  IVI U910 ( .A(n2522), .Z(n2118) );
  IVI U911 ( .A(n2073), .Z(speed[2]) );
  AN3 U912 ( .A(speed[2]), .B(speed[1]), .C(speed[3]), .Z(n1852) );
  IVI U913 ( .A(n2112), .Z(n2120) );
  ND2I U914 ( .A(n2191), .B(n2192), .Z(n2235) );
  INVX1 U915 ( .A(n2121), .Y(n2183) );
  NAND2X1 U916 ( .A(n2372), .B(n2371), .Y(n2121) );
  OR2X1 U917 ( .A(n2108), .B(n2143), .Y(n2371) );
  AN2I U918 ( .A(n2256), .B(n2257), .Z(n2122) );
  IVI U919 ( .A(n2155), .Z(n2123) );
  AN2I U920 ( .A(n2413), .B(n2444), .Z(n2124) );
  AN2I U921 ( .A(n2372), .B(n2158), .Z(n2125) );
  ND2I U922 ( .A(n2283), .B(n2282), .Z(n2127) );
  MUX21LP U923 ( .A(n845), .B(N46), .S(accel), .Z(n2303) );
  AO3P U924 ( .A(n2302), .B(n2069), .C(n2301), .D(n2300), .Z(n2368) );
  ND2I U925 ( .A(n2526), .B(n2525), .Z(n2128) );
  ND2I U926 ( .A(n2219), .B(n2145), .Z(n2129) );
  IVI U927 ( .A(n2122), .Z(n2130) );
  IVI U928 ( .A(n2130), .Z(n2131) );
  ND2I U929 ( .A(n2464), .B(n2463), .Z(n2132) );
  IVI U930 ( .A(n2139), .Z(n2133) );
  IVI U931 ( .A(n2133), .Z(n2134) );
  ND2I U932 ( .A(coast), .B(n2127), .Z(n2135) );
  OR2I U933 ( .A(n2266), .B(reset), .Z(n2136) );
  NR2I U934 ( .A(n2137), .B(reset), .Z(N259) );
  ND2I U935 ( .A(n2476), .B(n2475), .Z(n2138) );
  ND2I U936 ( .A(accel), .B(n2116), .Z(n2139) );
  AND2X1 U937 ( .A(n2369), .B(n2029), .Y(n2154) );
  OR2X1 U938 ( .A(n2154), .B(n2153), .Y(n2372) );
  IVI U939 ( .A(n2141), .Z(n2469) );
  AN2I U940 ( .A(n2411), .B(n2410), .Z(n2141) );
  ND2I U941 ( .A(n2181), .B(n2182), .Z(n2142) );
  B4IP U942 ( .A(n2432), .Z(n2143) );
  B4IP U943 ( .A(n2234), .Z(n2251) );
  NR2I U944 ( .A(n2625), .B(n2116), .Z(n2310) );
  AN2I U945 ( .A(n2390), .B(n2215), .Z(n2308) );
  AN2I U946 ( .A(n2568), .B(n2591), .Z(n2146) );
  IVI U947 ( .A(n2134), .Z(n2383) );
  IVI U948 ( .A(n2307), .Z(n2147) );
  NR2I U949 ( .A(n2149), .B(n2308), .Z(n2148) );
  ND2I U950 ( .A(n2309), .B(n2147), .Z(n2149) );
  IVI U951 ( .A(n2152), .Z(n2163) );
  B4IP U952 ( .A(n2288), .Z(n2031) );
  AN2I U953 ( .A(n2256), .B(n2257), .Z(n2150) );
  IVI U954 ( .A(n2129), .Z(n2151) );
  AN2I U955 ( .A(set), .B(n2159), .Z(n2152) );
  ND2I U956 ( .A(n2172), .B(n2146), .Z(n2494) );
  B4IP U957 ( .A(n2368), .Z(n2153) );
  B4IP U958 ( .A(n2573), .Z(n2258) );
  ND2I U959 ( .A(n2425), .B(n2424), .Z(n2155) );
  ND2I U960 ( .A(n2141), .B(n2247), .Z(n2156) );
  IVI U961 ( .A(n2527), .Z(n2157) );
  NR2I U962 ( .A(n2573), .B(n2164), .Z(n2429) );
  ND2I U963 ( .A(n2370), .B(n2432), .Z(n2158) );
  ND2I U964 ( .A(n2509), .B(n2508), .Z(n2159) );
  IVI U965 ( .A(n2430), .Z(n2160) );
  IVI U966 ( .A(n2139), .Z(n2161) );
  ND2I U967 ( .A(n2511), .B(n2656), .Z(n2162) );
  ND2I U968 ( .A(n2372), .B(n2158), .Z(n2164) );
  ND2I U969 ( .A(n2423), .B(n2422), .Z(n2165) );
  ND2I U970 ( .A(n2423), .B(n2422), .Z(n2166) );
  ND2I U971 ( .A(n2514), .B(n2117), .Z(n2167) );
  B2IP U972 ( .A(n2667), .Z2(n2168) );
  ND2I U973 ( .A(n2423), .B(n2422), .Z(n2581) );
  IVI U974 ( .A(n2285), .Z(n2667) );
  ND2I U975 ( .A(n2638), .B(brake), .Z(n2170) );
  ND2I U976 ( .A(n2170), .B(n2171), .Z(n179) );
  ND2I U977 ( .A(n2579), .B(n2493), .Z(n2172) );
  NAND2X1 U978 ( .A(n2175), .B(n2173), .Y(n2197) );
  AND2X1 U979 ( .A(n2176), .B(n2366), .Y(n2173) );
  NAND2X1 U980 ( .A(n2175), .B(n2174), .Y(n2198) );
  AND2X1 U981 ( .A(n2176), .B(n2070), .Y(n2174) );
  OR2X1 U982 ( .A(n2217), .B(n2216), .Y(n2175) );
  OR2X2 U983 ( .A(n2360), .B(n2030), .Y(n2176) );
  MUX21LP U984 ( .A(n2567), .B(n2373), .S(n2164), .Z(n2405) );
  MUX21LP U985 ( .A(n841), .B(N50), .S(accel), .Z(n2177) );
  NAND2X1 U986 ( .A(n2184), .B(n2242), .Y(n2178) );
  NAND2X1 U987 ( .A(n2395), .B(n2184), .Y(n2179) );
  NAND2X1 U988 ( .A(n2242), .B(n2395), .Y(n2180) );
  NAND3X1 U989 ( .A(n2178), .B(n2180), .C(n2179), .Y(n2396) );
  MUX21LP U990 ( .A(speed[3]), .B(N39), .S(n2121), .Z(n2453) );
  MUX21LP U991 ( .A(N37), .B(speed[1]), .S(n2183), .Z(n2255) );
  ND2I U992 ( .A(N36), .B(n2121), .Z(n2181) );
  ND2I U993 ( .A(speed[0]), .B(n2183), .Z(n2182) );
  AND2X1 U994 ( .A(n2394), .B(n2478), .Y(n2184) );
  ND2I U995 ( .A(n2058), .B(n2653), .Z(n2186) );
  ND2I U996 ( .A(n2186), .B(n2187), .Z(n2228) );
  OR2P U997 ( .A(brake), .B(n2658), .Z(n2187) );
  AN2I U998 ( .A(n2126), .B(n2659), .Z(n2188) );
  NOR2X1 U999 ( .A(n2051), .B(n2407), .Y(n2189) );
  INVX1 U1000 ( .A(n2220), .Y(n2190) );
  OR2X1 U1001 ( .A(n2190), .B(n2189), .Y(n2408) );
  ND2I U1002 ( .A(N40), .B(n2121), .Z(n2191) );
  ND2I U1003 ( .A(n838), .B(n2183), .Z(n2192) );
  ND2I U1004 ( .A(N38), .B(n2121), .Z(n2193) );
  ND2I U1005 ( .A(speed[2]), .B(n2183), .Z(n2194) );
  ND2I U1006 ( .A(n2193), .B(n2194), .Z(n2195) );
  ND2I U1007 ( .A(n2155), .B(n2659), .Z(n2196) );
  NAND2X1 U1008 ( .A(n2366), .B(n2070), .Y(n2199) );
  NAND3X1 U1009 ( .A(n2199), .B(n2197), .C(n2198), .Y(n2369) );
  NAND2X1 U1010 ( .A(n2252), .B(n2396), .Y(n2200) );
  NAND2X1 U1011 ( .A(n2252), .B(n2218), .Y(n2201) );
  NAND2X1 U1012 ( .A(n2218), .B(n2396), .Y(n2202) );
  NAND3X1 U1013 ( .A(n2201), .B(n2202), .C(n2200), .Y(n2399) );
  NAND2X1 U1014 ( .A(n2398), .B(n2062), .Y(n2203) );
  NAND2X1 U1015 ( .A(n2401), .B(n2402), .Y(n2204) );
  NAND3X1 U1016 ( .A(n2204), .B(n2203), .C(n2061), .Y(n2403) );
  NAND2X1 U1017 ( .A(n2353), .B(n2352), .Y(n2205) );
  NAND2X1 U1018 ( .A(n2213), .B(n2353), .Y(n2206) );
  NAND2X1 U1019 ( .A(n2352), .B(n2213), .Y(n2207) );
  NAND3X1 U1020 ( .A(n2207), .B(n2205), .C(n2206), .Y(n2360) );
  NAND2X1 U1021 ( .A(n2113), .B(n2254), .Y(n2208) );
  NAND2X1 U1022 ( .A(n2254), .B(n2404), .Y(n2209) );
  NAND3X1 U1023 ( .A(n2208), .B(n2209), .C(n2055), .Y(n2407) );
  NAND2X1 U1024 ( .A(n2210), .B(n2211), .Y(n2212) );
  B4IP U1025 ( .A(n2110), .Z(n2210) );
  INVX1 U1026 ( .A(n2403), .Y(n2211) );
  B4IP U1027 ( .A(n2255), .Z(n2248) );
  OR2I U1028 ( .A(n2132), .B(n2101), .Z(n2601) );
  AO3P U1029 ( .A(n2429), .B(n2428), .C(n2427), .D(n2426), .Z(n2430) );
  B4IP U1030 ( .A(n2381), .Z(n2400) );
  B4IP U1031 ( .A(n2144), .Z(n2478) );
  NOR2X1 U1032 ( .A(reset), .B(n2214), .Y(n2213) );
  B4IP U1033 ( .A(n838), .Z(n2214) );
  IVI U1034 ( .A(n2347), .Z(n2215) );
  INVX1 U1035 ( .A(n2290), .Y(n2030) );
  IVI U1036 ( .A(n2215), .Z(n2219) );
  B4IP U1037 ( .A(n2377), .Z(n2216) );
  B4IP U1038 ( .A(n2432), .Z(n2029) );
  AO3P U1039 ( .A(n1307), .B(N202), .C(N200), .D(N201), .Z(n2649) );
  B4IP U1040 ( .A(n2413), .Z(n2244) );
  B4IP U1041 ( .A(n2388), .Z(n2231) );
  B4IP U1042 ( .A(n2387), .Z(n2230) );
  AND2X1 U1043 ( .A(n2231), .B(n2230), .Y(n2218) );
  IVI U1044 ( .A(n2376), .Z(n2223) );
  OR2I U1045 ( .A(n2236), .B(n2237), .Z(n1738) );
  IVI U1046 ( .A(n2603), .Z(n2605) );
  IVI U1047 ( .A(n2455), .Z(n2412) );
  IVI U1048 ( .A(n2338), .Z(n2274) );
  AN2I U1049 ( .A(n2497), .B(n2496), .Z(n2221) );
  IVI U1050 ( .A(n2582), .Z(n2419) );
  IVI U1051 ( .A(n2598), .Z(n2602) );
  IVI U1052 ( .A(n2558), .Z(n2559) );
  IVI U1053 ( .A(n2550), .Z(n2551) );
  IVI U1054 ( .A(n2384), .Z(n2536) );
  IVI U1055 ( .A(n2647), .Z(n2638) );
  AN2I U1056 ( .A(n2120), .B(n2550), .Z(n2224) );
  IVI U1057 ( .A(n2378), .Z(n2512) );
  IVI U1058 ( .A(n2444), .Z(n2445) );
  IVI U1059 ( .A(n2484), .Z(n2314) );
  IVI U1060 ( .A(n2584), .Z(n2487) );
  AN2I U1061 ( .A(n2447), .B(n2498), .Z(n2225) );
  IVI U1062 ( .A(n2457), .Z(n2289) );
  AN2I U1063 ( .A(n2458), .B(n2457), .Z(n2226) );
  AN2I U1064 ( .A(n2333), .B(n2332), .Z(n2227) );
  B4IP U1065 ( .A(n2227), .Z(n2346) );
  IVI U1066 ( .A(n2336), .Z(n2272) );
  IVI U1067 ( .A(n2320), .Z(n2271) );
  IVI U1068 ( .A(n2468), .Z(n2411) );
  IVI U1069 ( .A(n2496), .Z(n2416) );
  IVI U1070 ( .A(n2128), .Z(n2648) );
  IVI U1071 ( .A(n2612), .Z(n2613) );
  IVI U1072 ( .A(n2297), .Z(n2354) );
  IVI U1073 ( .A(n2278), .Z(n2304) );
  AN2I U1074 ( .A(speed[6]), .B(n2518), .Z(n2367) );
  IVI U1075 ( .A(n2604), .Z(n2606) );
  IVI U1076 ( .A(n2643), .Z(n2644) );
  IVI U1077 ( .A(n2437), .Z(n2406) );
  IVI U1078 ( .A(N42), .Z(n2373) );
  ND2I U1079 ( .A(n2048), .B(n2233), .Z(n2232) );
  AN2I U1080 ( .A(n2392), .B(n2391), .Z(n2233) );
  IVI U1081 ( .A(n2319), .Z(n2321) );
  IVI U1082 ( .A(n2247), .Z(n2454) );
  MUX21L U1083 ( .A(N40), .B(n2597), .S(n2125), .Z(n2444) );
  IVI U1084 ( .A(n2303), .Z(n2625) );
  IVI U1085 ( .A(n2335), .Z(n2337) );
  AN2I U1086 ( .A(n2351), .B(n2350), .Z(n2234) );
  IVI U1087 ( .A(n2415), .Z(n2414) );
  NR2I U1088 ( .A(n2589), .B(n2588), .Z(n2645) );
  AO3 U1089 ( .A(n2029), .B(n2433), .C(n2428), .D(n2659), .Z(n2427) );
  IVI U1090 ( .A(n2582), .Z(n2583) );
  IVI U1091 ( .A(n2427), .Z(n2294) );
  IVI U1092 ( .A(n2498), .Z(n2291) );
  IVI U1093 ( .A(n2465), .Z(n2287) );
  IVI U1094 ( .A(n2499), .Z(n2293) );
  IVI U1095 ( .A(n2428), .Z(n2655) );
  IVI U1096 ( .A(n2609), .Z(n2506) );
  IVI U1097 ( .A(n2327), .Z(n2328) );
  MUX21L U1098 ( .A(n843), .B(N48), .S(accel), .Z(n2319) );
  MUX21L U1099 ( .A(N43), .B(speed[7]), .S(n2183), .Z(n2437) );
  MUX21L U1100 ( .A(cruise_speed[3]), .B(n2157), .S(accel), .Z(n2335) );
  MUX21L U1101 ( .A(n2640), .B(n2639), .S(brake), .Z(n2642) );
  ND2I U1102 ( .A(n2600), .B(n2599), .Z(n2236) );
  MUX21L U1103 ( .A(N42), .B(speed[6]), .S(n2125), .Z(n2415) );
  MUX21L U1104 ( .A(n2594), .B(n2593), .S(brake), .Z(n2596) );
  MUX21L U1105 ( .A(n2571), .B(n2570), .S(brake), .Z(n2577) );
  MUX21H U1106 ( .A(n2579), .B(n2172), .S(brake), .Z(n2238) );
  AN2I U1107 ( .A(n2575), .B(n2574), .Z(n2239) );
  IVI U1108 ( .A(reset), .Z(n2518) );
  AN2I U1109 ( .A(n2240), .B(n2241), .Z(n2660) );
  AN2I U1110 ( .A(n2567), .B(n2269), .Z(n2241) );
  MUX21H U1111 ( .A(speed[5]), .B(n2024), .S(n2660), .Z(n168) );
  MUX21H U1112 ( .A(speed[3]), .B(n2021), .S(n2660), .Z(n170) );
  MUX21H U1113 ( .A(speed[2]), .B(n2022), .S(n2660), .Z(n2665) );
  MUX21L U1114 ( .A(n2072), .B(n2089), .S(n2660), .Z(n2664) );
  MUX21H U1115 ( .A(speed[0]), .B(n2027), .S(n2660), .Z(n2661) );
  BUFX2 U1116 ( .A(n2248), .Y(n2242) );
  MUX21L U1117 ( .A(n2482), .B(n2481), .S(n2125), .Z(n2483) );
  MUX21L U1118 ( .A(N37), .B(speed[1]), .S(n2125), .Z(n2477) );
  INVX1 U1119 ( .A(n2114), .Y(n2243) );
  B4IP U1120 ( .A(n2235), .Z(n2245) );
  B4IP U1121 ( .A(n2453), .Z(n2246) );
  INVX1 U1122 ( .A(n2246), .Y(n2247) );
  B4IP U1123 ( .A(n1231), .Z(n2249) );
  INVX1 U1124 ( .A(n2249), .Y(n2250) );
  IVI U1125 ( .A(n2332), .Z(n1231) );
  INVX1 U1126 ( .A(n2245), .Y(n2401) );
  BUFX2 U1127 ( .A(n2467), .Y(n2252) );
  B4IP U1128 ( .A(n2410), .Z(n2467) );
  B4IP U1129 ( .A(n2405), .Z(n2253) );
  INVX1 U1130 ( .A(n2253), .Y(n2254) );
  ND2I U1131 ( .A(n2159), .B(set), .Z(n2256) );
  AN2I U1132 ( .A(n2256), .B(n2257), .Z(n2628) );
  AN2I U1133 ( .A(n2521), .B(n2518), .Z(n2257) );
  ND2I U1134 ( .A(n2258), .B(n2259), .Z(n2423) );
  NR2I U1135 ( .A(n2428), .B(n2125), .Z(n2259) );
  IVI U1136 ( .A(n2136), .Z(n2260) );
  IVI U1137 ( .A(n2640), .Z(n2443) );
  IVI U1138 ( .A(n2264), .Z(N267) );
  NAND2X1 U1139 ( .A(n2573), .B(n2520), .Y(n2582) );
  OR2I U1140 ( .A(n2265), .B(reset), .Z(n2264) );
  OR2I U1141 ( .A(n2262), .B(reset), .Z(n2261) );
  IVI U1142 ( .A(n2261), .Z(n2263) );
  IVI U1143 ( .A(n2519), .Z(n2389) );
  IVI U1144 ( .A(n2393), .Z(n2394) );
  IVI U1145 ( .A(n2334), .Z(n2333) );
  B4IP U1146 ( .A(n2267), .Z(n2345) );
  B4IP U1147 ( .A(n2286), .Z(n2668) );
  NAND2X1 U1148 ( .A(n2409), .B(n2408), .Y(n2573) );
  NAND2X1 U1149 ( .A(n2051), .B(n2057), .Y(n2409) );
  OR2P U1150 ( .A(n2268), .B(reset), .Z(n2292) );
  IVI U1151 ( .A(n2362), .Z(n2299) );
  INVX1 U1152 ( .A(n2049), .Y(n2366) );
  B4IP U1153 ( .A(n2292), .Z(n1474) );
  AND2X1 U1154 ( .A(n2345), .B(n2346), .Y(n2353) );
  NAND2X1 U1155 ( .A(n2247), .B(n2397), .Y(n2398) );
  INVX1 U1156 ( .A(n2251), .Y(n2352) );
  MUX21L U1157 ( .A(n2028), .B(n2090), .S(n2660), .Z(n169) );
  IVI U1158 ( .A(n2430), .Z(n2633) );
  IVI U1159 ( .A(n2571), .Z(n2476) );
  NAND2X1 U1160 ( .A(n2400), .B(n2399), .Y(n2397) );
  IVI U1161 ( .A(n2355), .Z(n2298) );
  IVI U1162 ( .A(n2594), .Z(n2464) );
  IVI U1163 ( .A(n2492), .Z(n2579) );
  IVI U1164 ( .A(speed[6]), .Z(n2567) );
  IVI U1165 ( .A(n2028), .Z(n2597) );
  ND2I U1166 ( .A(n2660), .B(n2026), .Z(n2270) );
  ND2I U1167 ( .A(n2240), .B(n2270), .Z(n166) );
  NR2I U1168 ( .A(n159), .B(reset), .Z(N255) );
  AN2I U1169 ( .A(n839), .B(n2518), .Z(N257) );
  NR2I U1170 ( .A(n2019), .B(reset), .Z(N261) );
  ND2I U1171 ( .A(speed[7]), .B(n2518), .Z(n2432) );
  ND2I U1172 ( .A(speed[5]), .B(n2518), .Z(n2290) );
  ND2I U1173 ( .A(n2597), .B(n2518), .Z(n2288) );
  ND2I U1174 ( .A(speed[3]), .B(n2518), .Z(n2332) );
  ND2I U1175 ( .A(n2669), .B(n2518), .Z(n2286) );
  ND2I U1176 ( .A(speed[1]), .B(n2518), .Z(n2285) );
  ND2I U1177 ( .A(speed[0]), .B(n2518), .Z(n2585) );
  IVAP U1178 ( .A(n2585), .Z(n2032) );
  ND2I U1179 ( .A(n2303), .B(n2278), .Z(n2320) );
  ND2I U1180 ( .A(n2271), .B(n2319), .Z(n2336) );
  ND2I U1181 ( .A(n2272), .B(n2335), .Z(n2338) );
  IVI U1182 ( .A(N50), .Z(n2515) );
  ND2I U1183 ( .A(n2338), .B(n2273), .Z(n2275) );
  ND2I U1184 ( .A(n2274), .B(n2177), .Z(n2355) );
  ND2I U1185 ( .A(n2275), .B(n2355), .Z(n2378) );
  MUX21LP U1186 ( .A(cruise_speed[6]), .B(N52), .S(accel), .Z(n2361) );
  MUX21LP U1187 ( .A(cruise_speed[7]), .B(N53), .S(accel), .Z(n2614) );
  AN2I U1188 ( .A(n2361), .B(n2614), .Z(n2283) );
  ND2I U1189 ( .A(n843), .B(cruise_speed[3]), .Z(n2277) );
  ND2I U1190 ( .A(N49), .B(N48), .Z(n2276) );
  ND2I U1191 ( .A(n2279), .B(n2304), .Z(n2280) );
  ND2I U1192 ( .A(n2177), .B(n2280), .Z(n2281) );
  ND2I U1193 ( .A(n2281), .B(n2354), .Z(n2282) );
  ND2I U1194 ( .A(n2283), .B(n2282), .Z(n2284) );
  ND2I U1195 ( .A(coast), .B(n2284), .Z(n2347) );
  ND2I U1196 ( .A(cruise_on), .B(n2518), .Z(n2428) );
  IVI U1197 ( .A(throttle), .Z(n2422) );
  ND2I U1198 ( .A(n2655), .B(n2422), .Z(n2572) );
  NR2I U1199 ( .A(n2219), .B(n2572), .Z(n2511) );
  ND2I U1200 ( .A(n2585), .B(n2285), .Z(n2484) );
  ND2I U1201 ( .A(n2314), .B(n2286), .Z(n2465) );
  ND2I U1202 ( .A(n2287), .B(n2332), .Z(n2457) );
  ND2I U1203 ( .A(n2289), .B(n2288), .Z(n2498) );
  ND2I U1204 ( .A(n2291), .B(n2290), .Z(n2499) );
  ND2I U1205 ( .A(n2293), .B(n2292), .Z(n2433) );
  IVI U1206 ( .A(brake), .Z(n2659) );
  ND2I U1207 ( .A(n2294), .B(n2422), .Z(n2584) );
  ND2I U1208 ( .A(n1474), .B(n2499), .Z(n2295) );
  ND2I U1209 ( .A(n2295), .B(n2433), .Z(n2296) );
  ND2I U1210 ( .A(n2487), .B(n2296), .Z(n2421) );
  IVAP U1211 ( .A(n2572), .Z(n2520) );
  ND2I U1212 ( .A(n2298), .B(n2044), .Z(n2362) );
  ND2I U1213 ( .A(n2299), .B(n2043), .Z(n2612) );
  ND2I U1214 ( .A(n2120), .B(n2612), .Z(n2302) );
  ND2I U1215 ( .A(accel), .B(n2135), .Z(n2513) );
  ND2I U1216 ( .A(n2083), .B(n2161), .Z(n2301) );
  ND2I U1217 ( .A(n2112), .B(n2145), .Z(n2519) );
  ND2I U1218 ( .A(n2389), .B(cruise_speed[7]), .Z(n2300) );
  ND2I U1219 ( .A(n2625), .B(n2304), .Z(n2305) );
  ND2I U1220 ( .A(n2305), .B(n2320), .Z(n2390) );
  IVI U1221 ( .A(n844), .Z(n2306) );
  NR2I U1222 ( .A(n2519), .B(n2306), .Z(n2307) );
  ND2I U1223 ( .A(n2047), .B(n2161), .Z(n2309) );
  NR2I U1224 ( .A(n2263), .B(n2513), .Z(n2311) );
  NR2I U1225 ( .A(n2311), .B(n2310), .Z(n2313) );
  ND2I U1226 ( .A(n845), .B(n2389), .Z(n2312) );
  ND2I U1227 ( .A(n2313), .B(n2312), .Z(n2393) );
  ND2I U1228 ( .A(n2314), .B(n2393), .Z(n2315) );
  ND2I U1229 ( .A(n2148), .B(n2315), .Z(n2318) );
  ND2I U1230 ( .A(n2393), .B(n2585), .Z(n2316) );
  ND2I U1231 ( .A(n2667), .B(n2316), .Z(n2317) );
  ND2I U1232 ( .A(n2318), .B(n2317), .Z(n2329) );
  ND2I U1233 ( .A(n2668), .B(n2329), .Z(n2331) );
  ND2I U1234 ( .A(n2321), .B(n2320), .Z(n2322) );
  ND2I U1235 ( .A(n2322), .B(n2336), .Z(n2384) );
  NR2I U1236 ( .A(n2536), .B(n2219), .Z(n2324) );
  IVI U1237 ( .A(N48), .Z(n2535) );
  NR2I U1238 ( .A(n2535), .B(n2134), .Z(n2323) );
  NR2I U1239 ( .A(n2324), .B(n2323), .Z(n2326) );
  ND2I U1240 ( .A(n2389), .B(n843), .Z(n2325) );
  ND2I U1241 ( .A(n2326), .B(n2325), .Z(n2327) );
  AO7P U1242 ( .A(n2668), .B(n2329), .C(n2328), .Z(n2330) );
  ND2I U1243 ( .A(n2331), .B(n2330), .Z(n2334) );
  ND2I U1244 ( .A(n2250), .B(n2334), .Z(n2344) );
  ND2I U1245 ( .A(n2337), .B(n2336), .Z(n2339) );
  AN2I U1246 ( .A(n2339), .B(n2338), .Z(n2528) );
  NR2I U1247 ( .A(n2528), .B(n2219), .Z(n2341) );
  NR2I U1248 ( .A(n2086), .B(n2129), .Z(n2340) );
  NR2I U1249 ( .A(n2341), .B(n2340), .Z(n2343) );
  ND2I U1250 ( .A(n2383), .B(n2157), .Z(n2342) );
  ND2I U1251 ( .A(n2343), .B(n2342), .Z(n2381) );
  NR2I U1252 ( .A(n2512), .B(n2219), .Z(n2349) );
  NR2I U1253 ( .A(n2118), .B(n2129), .Z(n2348) );
  NR2I U1254 ( .A(n2349), .B(n2348), .Z(n2351) );
  ND2I U1255 ( .A(n2383), .B(N50), .Z(n2350) );
  ND2I U1256 ( .A(n2355), .B(n2045), .Z(n2356) );
  ND2I U1257 ( .A(n2356), .B(n2362), .Z(n2550) );
  IVI U1258 ( .A(N51), .Z(n2549) );
  NR2I U1259 ( .A(n2109), .B(n2549), .Z(n2357) );
  NR2I U1260 ( .A(n2224), .B(n2357), .Z(n2359) );
  ND2I U1261 ( .A(n840), .B(n2389), .Z(n2358) );
  ND2I U1262 ( .A(n2085), .B(n2383), .Z(n2375) );
  ND2I U1263 ( .A(n2362), .B(n2042), .Z(n2363) );
  ND2I U1264 ( .A(n2363), .B(n2612), .Z(n2558) );
  ND2I U1265 ( .A(n2120), .B(n2558), .Z(n2374) );
  ND2I U1266 ( .A(cruise_speed[6]), .B(n2151), .Z(n2364) );
  ND2I U1267 ( .A(n2223), .B(n2364), .Z(n2365) );
  ND2I U1268 ( .A(n2375), .B(n2374), .Z(n2376) );
  IVI U1269 ( .A(n2019), .Z(n2522) );
  ND2I U1270 ( .A(n2151), .B(n2522), .Z(n2380) );
  ND2I U1271 ( .A(n2120), .B(n2378), .Z(n2379) );
  IVI U1272 ( .A(n843), .Z(n2382) );
  NR2I U1273 ( .A(n2382), .B(n2129), .Z(n2388) );
  ND2I U1274 ( .A(n2383), .B(N48), .Z(n2386) );
  ND2I U1275 ( .A(n2120), .B(n2384), .Z(n2385) );
  ND2I U1276 ( .A(n2386), .B(n2385), .Z(n2387) );
  ND2I U1277 ( .A(n844), .B(n2151), .Z(n2392) );
  ND2I U1278 ( .A(n2120), .B(n2390), .Z(n2391) );
  IVI U1279 ( .A(N37), .Z(n2480) );
  ND2I U1280 ( .A(n2053), .B(n2477), .Z(n2468) );
  ND2I U1281 ( .A(n2141), .B(n2247), .Z(n2455) );
  ND2I U1282 ( .A(n2412), .B(n2444), .Z(n2495) );
  ND2I U1283 ( .A(n2124), .B(n2412), .Z(n2496) );
  ND2I U1284 ( .A(n2496), .B(n2414), .Z(n2417) );
  ND2I U1285 ( .A(n2416), .B(n2415), .Z(n2438) );
  ND2I U1286 ( .A(n2417), .B(n2438), .Z(n2418) );
  ND2I U1287 ( .A(n2419), .B(n2418), .Z(n2420) );
  AN2I U1288 ( .A(n2421), .B(n2420), .Z(n2425) );
  ND2I U1289 ( .A(N42), .B(n2165), .Z(n2424) );
  NR2I U1290 ( .A(throttle), .B(reset), .Z(n2426) );
  ND2I U1291 ( .A(n2160), .B(speed[6]), .Z(n2431) );
  ND2I U1292 ( .A(n2123), .B(n2431), .Z(n2637) );
  ND2I U1293 ( .A(N43), .B(n2165), .Z(n2436) );
  NR2I U1294 ( .A(n2584), .B(n2432), .Z(n2434) );
  ND2I U1295 ( .A(n2434), .B(n2433), .Z(n2435) );
  AN2I U1296 ( .A(n2436), .B(n2435), .Z(n2441) );
  NR2I U1297 ( .A(n2437), .B(n2582), .Z(n2439) );
  ND2I U1298 ( .A(n2439), .B(n2438), .Z(n2440) );
  ND2I U1299 ( .A(n2441), .B(n2440), .Z(n2640) );
  ND2I U1300 ( .A(n2160), .B(speed[7]), .Z(n2442) );
  ND2I U1301 ( .A(n2443), .B(n2442), .Z(n2643) );
  NR2I U1302 ( .A(n2637), .B(n2643), .Z(n2509) );
  ND2I U1303 ( .A(n2445), .B(n2156), .Z(n2446) );
  NR2I U1304 ( .A(n2054), .B(n2582), .Z(n2449) );
  ND2I U1305 ( .A(n2031), .B(n2457), .Z(n2447) );
  NR2I U1306 ( .A(n2225), .B(n2584), .Z(n2448) );
  NR2I U1307 ( .A(n2449), .B(n2448), .Z(n2451) );
  ND2I U1308 ( .A(N40), .B(n2166), .Z(n2450) );
  ND2I U1309 ( .A(n2160), .B(n2597), .Z(n2452) );
  ND2I U1310 ( .A(n2064), .B(n2452), .Z(n2598) );
  ND2I U1311 ( .A(n2469), .B(n2454), .Z(n2456) );
  NR2I U1312 ( .A(n2075), .B(n2582), .Z(n2460) );
  ND2I U1313 ( .A(n2250), .B(n2465), .Z(n2458) );
  NR2I U1314 ( .A(n2226), .B(n2584), .Z(n2459) );
  NR2I U1315 ( .A(n2460), .B(n2459), .Z(n2462) );
  ND2I U1316 ( .A(N39), .B(n2581), .Z(n2461) );
  ND2I U1317 ( .A(n2462), .B(n2461), .Z(n2594) );
  ND2I U1318 ( .A(n2633), .B(speed[3]), .Z(n2463) );
  ND2I U1319 ( .A(n2464), .B(n2463), .Z(n2591) );
  ND2I U1320 ( .A(n2668), .B(n2484), .Z(n2466) );
  NR2I U1321 ( .A(n2088), .B(n2584), .Z(n2472) );
  ND2I U1322 ( .A(n2468), .B(n2252), .Z(n2470) );
  NR2I U1323 ( .A(n2076), .B(n2582), .Z(n2471) );
  NR2I U1324 ( .A(n2472), .B(n2471), .Z(n2474) );
  ND2I U1325 ( .A(N38), .B(n2581), .Z(n2473) );
  ND2I U1326 ( .A(n2474), .B(n2473), .Z(n2571) );
  ND2I U1327 ( .A(n2633), .B(speed[2]), .Z(n2475) );
  ND2I U1328 ( .A(n2476), .B(n2475), .Z(n2568) );
  ND2I U1329 ( .A(n2052), .B(n2477), .Z(n2479) );
  NR2I U1330 ( .A(N36), .B(n2480), .Z(n2482) );
  NR2I U1331 ( .A(speed[0]), .B(n2072), .Z(n2481) );
  ND2I U1332 ( .A(n2032), .B(n2168), .Z(n2485) );
  ND2I U1333 ( .A(n2485), .B(n2484), .Z(n2486) );
  ND2I U1334 ( .A(n2487), .B(n2486), .Z(n2488) );
  AN2I U1335 ( .A(n2489), .B(n2488), .Z(n2491) );
  ND2I U1336 ( .A(N37), .B(n2166), .Z(n2490) );
  ND2I U1337 ( .A(n2491), .B(n2490), .Z(n2492) );
  ND2I U1338 ( .A(n2160), .B(speed[1]), .Z(n2493) );
  ND2I U1339 ( .A(n2579), .B(n2493), .Z(n2578) );
  ND2I U1340 ( .A(n2602), .B(n2494), .Z(n2507) );
  ND2I U1341 ( .A(n2495), .B(n2244), .Z(n2497) );
  NR2I U1342 ( .A(n2221), .B(n2582), .Z(n2502) );
  ND2I U1343 ( .A(n2030), .B(n2498), .Z(n2500) );
  NR2I U1344 ( .A(n2087), .B(n2584), .Z(n2501) );
  NR2I U1345 ( .A(n2502), .B(n2501), .Z(n2504) );
  ND2I U1346 ( .A(N41), .B(n2166), .Z(n2503) );
  ND2I U1347 ( .A(n2504), .B(n2503), .Z(n2609) );
  ND2I U1348 ( .A(n2160), .B(speed[5]), .Z(n2505) );
  ND2I U1349 ( .A(n2506), .B(n2505), .Z(n2604) );
  ND2I U1350 ( .A(n2507), .B(n2604), .Z(n2508) );
  ND2I U1351 ( .A(n2509), .B(n2508), .Z(n2510) );
  ND2I U1352 ( .A(set), .B(n2510), .Z(n2656) );
  ND2I U1353 ( .A(n2511), .B(n2656), .Z(n2624) );
  NR2I U1354 ( .A(n2512), .B(n2162), .Z(n2517) );
  NR2I U1355 ( .A(n2109), .B(n2572), .Z(n2514) );
  ND2I U1356 ( .A(n2514), .B(n2117), .Z(n2623) );
  NR2I U1357 ( .A(n2515), .B(n2095), .Z(n2516) );
  NR2I U1358 ( .A(n2517), .B(n2516), .Z(n2526) );
  ND2I U1359 ( .A(n2020), .B(n2152), .Z(n2524) );
  ND2I U1360 ( .A(n2520), .B(n2129), .Z(n2521) );
  ND2I U1361 ( .A(n2628), .B(n2522), .Z(n2523) );
  AN2I U1362 ( .A(n2524), .B(n2523), .Z(n2525) );
  IVI U1363 ( .A(N49), .Z(n2527) );
  NR2I U1364 ( .A(n2527), .B(n2167), .Z(n2530) );
  NR2I U1365 ( .A(n2528), .B(n2162), .Z(n2529) );
  NR2I U1366 ( .A(n2530), .B(n2529), .Z(n2534) );
  ND2I U1367 ( .A(n2021), .B(n2152), .Z(n2532) );
  ND2I U1368 ( .A(n2150), .B(cruise_speed[3]), .Z(n2531) );
  AN2I U1369 ( .A(n2532), .B(n2531), .Z(n2533) );
  ND2I U1370 ( .A(n2534), .B(n2533), .Z(N200) );
  NR2I U1371 ( .A(n2535), .B(n2167), .Z(n2538) );
  NR2I U1372 ( .A(n2536), .B(n2624), .Z(n2537) );
  NR2I U1373 ( .A(n2538), .B(n2537), .Z(n2542) );
  ND2I U1374 ( .A(n2022), .B(n2152), .Z(n2540) );
  ND2I U1375 ( .A(n2628), .B(n843), .Z(n2539) );
  AN2I U1376 ( .A(n2540), .B(n2539), .Z(n2541) );
  ND2I U1377 ( .A(n2542), .B(n2541), .Z(N201) );
  NR2I U1378 ( .A(n2077), .B(n2100), .Z(n2544) );
  NR2I U1379 ( .A(n2046), .B(n2095), .Z(n2543) );
  NR2I U1380 ( .A(n2544), .B(n2543), .Z(n2548) );
  ND2I U1381 ( .A(n2023), .B(n2152), .Z(n2546) );
  ND2I U1382 ( .A(n2150), .B(n844), .Z(n2545) );
  AN2I U1383 ( .A(n2546), .B(n2545), .Z(n2547) );
  ND2I U1384 ( .A(n2548), .B(n2547), .Z(N202) );
  NR2I U1385 ( .A(n2549), .B(n2167), .Z(n2553) );
  NR2I U1386 ( .A(n2551), .B(n2162), .Z(n2552) );
  NR2I U1387 ( .A(n2553), .B(n2552), .Z(n2557) );
  ND2I U1388 ( .A(n2024), .B(n2152), .Z(n2555) );
  ND2I U1389 ( .A(n2131), .B(n840), .Z(n2554) );
  AN2I U1390 ( .A(n2555), .B(n2554), .Z(n2556) );
  ND2I U1391 ( .A(n2557), .B(n2556), .Z(N198) );
  NR2I U1392 ( .A(n2084), .B(n2623), .Z(n2561) );
  NR2I U1393 ( .A(n2559), .B(n2100), .Z(n2560) );
  NR2I U1394 ( .A(n2561), .B(n2560), .Z(n2565) );
  ND2I U1395 ( .A(n2025), .B(n2152), .Z(n2563) );
  ND2I U1396 ( .A(n2115), .B(cruise_speed[6]), .Z(n2562) );
  AN2I U1397 ( .A(n2563), .B(n2562), .Z(n2564) );
  ND2I U1398 ( .A(n2565), .B(n2564), .Z(N197) );
  ND2I U1399 ( .A(n2660), .B(n2025), .Z(n2566) );
  ND2I U1400 ( .A(n2567), .B(n2566), .Z(n2666) );
  ND2I U1401 ( .A(n2578), .B(n2138), .Z(n2569) );
  ND2I U1402 ( .A(n2569), .B(n2101), .Z(n2570) );
  NR2I U1403 ( .A(n2572), .B(n2164), .Z(n2575) );
  NR2I U1404 ( .A(brake), .B(n2573), .Z(n2574) );
  ND2I U1405 ( .A(n2239), .B(speed[2]), .Z(n2576) );
  ND2I U1406 ( .A(n2577), .B(n2576), .Z(n1311) );
  ND2I U1407 ( .A(n2239), .B(speed[1]), .Z(n2580) );
  ND2I U1408 ( .A(n2580), .B(n2238), .Z(n174) );
  AN2I U1409 ( .A(N36), .B(n2165), .Z(n2589) );
  ND2I U1410 ( .A(n2583), .B(n2053), .Z(n2587) );
  ND2I U1411 ( .A(n2487), .B(n2585), .Z(n2586) );
  ND2I U1412 ( .A(n2587), .B(n2586), .Z(n2588) );
  ND2I U1413 ( .A(n2160), .B(speed[0]), .Z(n2590) );
  ND2I U1414 ( .A(n2645), .B(n2590), .Z(n2663) );
  ND2I U1415 ( .A(n2102), .B(n2132), .Z(n2592) );
  ND2I U1416 ( .A(n2592), .B(n2601), .Z(n2593) );
  ND2I U1417 ( .A(n2239), .B(speed[3]), .Z(n2595) );
  ND2I U1418 ( .A(n2596), .B(n2595), .Z(n176) );
  ND2I U1419 ( .A(n2239), .B(n2597), .Z(n2600) );
  ND2I U1420 ( .A(n2601), .B(n2598), .Z(n2599) );
  ND2I U1421 ( .A(n2105), .B(n2602), .Z(n2603) );
  ND2I U1422 ( .A(n2097), .B(n2604), .Z(n2607) );
  ND2I U1423 ( .A(n2606), .B(n2605), .Z(n2636) );
  ND2I U1424 ( .A(n2607), .B(n2636), .Z(n2608) );
  ND2I U1425 ( .A(n2239), .B(speed[5]), .Z(n2610) );
  ND2I U1426 ( .A(n2611), .B(n2610), .Z(n178) );
  ND2I U1427 ( .A(n2131), .B(cruise_speed[7]), .Z(n2617) );
  NR2I U1428 ( .A(n2613), .B(n2100), .Z(n2615) );
  ND2I U1429 ( .A(n2615), .B(n2068), .Z(n2616) );
  AN2I U1430 ( .A(n2617), .B(n2616), .Z(n2621) );
  NR2I U1431 ( .A(n2163), .B(n2091), .Z(n2619) );
  NR2I U1432 ( .A(n2082), .B(n2095), .Z(n2618) );
  NR2I U1433 ( .A(n2619), .B(n2618), .Z(n2620) );
  ND2I U1434 ( .A(n2621), .B(n2620), .Z(n2662) );
  IVI U1435 ( .A(N46), .Z(n2622) );
  NR2I U1436 ( .A(n2623), .B(n2622), .Z(n2627) );
  NR2I U1437 ( .A(n2625), .B(n2624), .Z(n2626) );
  NR2I U1438 ( .A(n2627), .B(n2626), .Z(n2632) );
  ND2I U1439 ( .A(n2027), .B(n2152), .Z(n2630) );
  ND2I U1440 ( .A(n2122), .B(n845), .Z(n2629) );
  AN2I U1441 ( .A(n2630), .B(n2629), .Z(n2631) );
  ND2I U1442 ( .A(n2632), .B(n2631), .Z(n1307) );
  ND2I U1443 ( .A(n2239), .B(speed[6]), .Z(n2635) );
  ND2I U1444 ( .A(n2123), .B(n2431), .Z(n2634) );
  ND2I U1445 ( .A(n2239), .B(speed[7]), .Z(n2641) );
  ND2I U1446 ( .A(n2642), .B(n2641), .Z(n180) );
  ND2I U1447 ( .A(n2645), .B(n2644), .Z(n2646) );
  NR2I U1448 ( .A(n2662), .B(N197), .Z(n2652) );
  ND2I U1449 ( .A(n2649), .B(n2648), .Z(n2650) );
  ND2I U1450 ( .A(n2650), .B(N198), .Z(n2651) );
  ND2I U1451 ( .A(n2652), .B(n2651), .Z(n2653) );
  IVI U1452 ( .A(cancel), .Z(n2654) );
  ND2I U1453 ( .A(n2655), .B(n2654), .Z(n2657) );
  AN2I U1454 ( .A(n2657), .B(n2163), .Z(n2658) );
endmodule

